* HW1 subcircuit John Sommers
.subckt SubCircuitHW1 in out gnd
R1 in out 1M
R2 out gnd 2M
.ends


